module sigmoid(clk,x,y);
input [15:0]x;
input clk;
output reg[15:0]y;
always @(posedge clk)
begin
if(x<16'b1111101000000000)begin//if x<-6, then y=0.
y=16'b0000000000000000;
end
//below is 'for a range of x, given a certain value to y'
else if(x<16'b1111101011100110)begin
y=16'b0000000000000001;
end
else if(x<16'b1111101101100110)begin
y=16'b0000000000000010;
end
else if(x<16'b1111101111001101)begin
y=16'b0000000000000011;
end
else if(x<16'b1111110000000000)begin
y=16'b0000000000000100;
end
else if(x<16'b1111110000110011)begin
y=16'b0000000000000101;
end
else if(x<16'b1111110001100110)begin
y=16'b0000000000000110;
end
else if(x<16'b1111110010000000)begin
y=16'b0000000000000111;
end
else if(x<16'b1111110010110011)begin
y=16'b0000000000001000;
end
else if(x<16'b1111110011001101)begin
y=16'b0000000000001001;
end
else if(x<16'b1111110011100110)begin
y=16'b0000000000001010;
end
else if(x<16'b1111110100000000)begin
y=16'b0000000000001011;
end
else if(x<16'b1111110100011010)begin
y=16'b0000000000001100;
end
else if(x<16'b1111110100110011)begin
y=16'b0000000000001101;
end
else if(x<16'b1111110101001101)begin
y=16'b0000000000001111;
end
else if(x<16'b1111110101100110)begin
y=16'b0000000000010000;
end
else if(x<16'b1111110110000000)begin
y=16'b0000000000010010;
end
else if(x<16'b1111110110011010)begin
y=16'b0000000000010011;
end
else if(x<16'b1111110110110011)begin
y=16'b0000000000010101;
end
else if(x<16'b1111110111001101)begin
y=16'b0000000000010111;
end
else if(x<16'b1111110111100110)begin
y=16'b0000000000011010;
end
else if(x<16'b1111111000000000)begin
y=16'b0000000000011100;
end
else if(x<16'b1111111000011010)begin
y=16'b0000000000011111;
end
else if(x<16'b1111111000110011)begin
y=16'b0000000000100001;
end
else if(x<16'b1111111001001101)begin
y=16'b0000000000100100;
end
else if(x<16'b1111111001100110)begin
y=16'b0000000000101000;
end
else if(x<16'b1111111010000000)begin
y=16'b0000000000101011;
end
else if(x<16'b1111111010011010)begin
y=16'b0000000000101111;
end
else if(x<16'b1111111010110011)begin
y=16'b0000000000110011;
end
else if(x<16'b1111111011001101)begin
y=16'b0000000000110111;
end
else if(x<16'b1111111011100110)begin
y=16'b0000000000111011;
end
else if(x<16'b1111111100000000)begin
y=16'b0000000001000000;
end
else if(x<16'b1111111100011010)begin
y=16'b0000000001000101;
end
else if(x<16'b1111111100110011)begin
y=16'b0000000001001010;
end
else if(x<16'b1111111101001101)begin
y=16'b0000000001001111;
end
else if(x<16'b1111111101100110)begin
y=16'b0000000001010101;
end
else if(x<16'b1111111110000000)begin
y=16'b0000000001011011;
end
else if(x<16'b1111111110011010)begin
y=16'b0000000001100001;
end
else if(x<16'b1111111110110011)begin
y=16'b0000000001100111;
end
else if(x<16'b1111111111001101)begin
y=16'b0000000001101101;
end
else if(x<16'b1111111111100110)begin
y=16'b0000000001110011;
end
else if(x<16'b0000000000000000)begin
y=16'b0000000001111010;
end
else if(x<16'b0000000000011010)begin
y=16'b0000000010000000;
end
else if(x<16'b0000000000110011)begin
y=16'b0000000010000110;
end
else if(x<16'b0000000001001101)begin
y=16'b0000000010001101;
end
else if(x<16'b0000000001100110)begin
y=16'b0000000010010011;
end
else if(x<16'b0000000010000000)begin
y=16'b0000000010011001;
end
else if(x<16'b0000000010011010)begin
y=16'b0000000010011111;
end
else if(x<16'b0000000010110011)begin
y=16'b0000000010100101;
end
else if(x<16'b0000000011001101)begin
y=16'b0000000010101011;
end
else if(x<16'b0000000011100110)begin
y=16'b0000000010110001;
end
else if(x<16'b0000000100000000)begin
y=16'b0000000010110110;
end
else if(x<16'b0000000100011010)begin
y=16'b0000000010111011;
end
else if(x<16'b0000000100110011)begin
y=16'b0000000011000000;
end
else if(x<16'b0000000101001101)begin
y=16'b0000000011000101;
end
else if(x<16'b0000000101100110)begin
y=16'b0000000011001001;
end
else if(x<16'b0000000110000000)begin
y=16'b0000000011001101;
end
else if(x<16'b0000000110011010)begin
y=16'b0000000011010001;
end
else if(x<16'b0000000110110011)begin
y=16'b0000000011010101;
end
else if(x<16'b0000000111001101)begin
y=16'b0000000011011000;
end
else if(x<16'b0000000111100110)begin
y=16'b0000000011011100;
end
else if(x<16'b0000001000000000)begin
y=16'b0000000011011111;
end
else if(x<16'b0000001000011010)begin
y=16'b0000000011100001;
end
else if(x<16'b0000001000110011)begin
y=16'b0000000011100100;
end
else if(x<16'b0000001001001101)begin
y=16'b0000000011100110;
end
else if(x<16'b0000001001100110)begin
y=16'b0000000011101001;
end
else if(x<16'b0000001010000000)begin
y=16'b0000000011101011;
end
else if(x<16'b0000001010011010)begin
y=16'b0000000011101101;
end
else if(x<16'b0000001010110011)begin
y=16'b0000000011101110;
end
else if(x<16'b0000001011001101)begin
y=16'b0000000011110000;
end
else if(x<16'b0000001011100110)begin
y=16'b0000000011110001;
end
else if(x<16'b0000001100000000)begin
y=16'b0000000011110011;
end
else if(x<16'b0000001100011010)begin
y=16'b0000000011110100;
end
else if(x<16'b0000001100110011)begin
y=16'b0000000011110101;
end
else if(x<16'b0000001101001101)begin
y=16'b0000000011110110;
end
else if(x<16'b0000001101100110)begin
y=16'b0000000011110111;
end
else if(x<16'b0000001110011010)begin
y=16'b0000000011111000;
end
else if(x<16'b0000001110110011)begin
y=16'b0000000011111001;
end
else if(x<16'b0000001111100110)begin
y=16'b0000000011111010;
end
else if(x<16'b0000010000011010)begin
y=16'b0000000011111011;
end
else if(x<16'b0000010001001101)begin
y=16'b0000000011111100;
end
else if(x<16'b0000010010110011)begin
y=16'b0000000011111101;
end
else if(x<16'b0000010100110011)begin
y=16'b0000000011111110;
end
else if(x<=16'b0000011000000000)begin
y=16'b0000000011111111;
end
else begin// if x>6,then y=1.
y=16'b0000000100000000;
end
end//end always
endmodule


